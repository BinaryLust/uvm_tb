
package div_pkg;

    import uvm_pkg::*;
	
    `include "div_random_item.svh"
	`include "div_constrained_random_item.svh"
	`include "div_output_trans.svh"
	
	`include "div_driver.svh"
	`include "div_input_monitor.svh"
	`include "div_output_monitor.svh"
	`include "div_sequencer.svh"
	`include "random_sequence.svh"
	`include "div_agent.svh"
	`include "div_coverage.svh"
	`include "div_scoreboard.svh"
	`include "div_env.svh"
	`include "base_test.svh"
	
endpackage

