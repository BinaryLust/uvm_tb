

`include "uvm_macros.svh"

module dut(dut_if dif);
    /*import uvm_pkg::*;
	always @(posedge dif.clk) begin
	    if(!dif.reset) begin
		    `uvm_info("DUT", $sformatf("opA = %h, opB = %h", dif.opA, dif.opB), UVM_MEDIUM)
		end
	end*/
endmodule

